module user_project_wrapper(
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif
    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);
	assign wbs_ack_o = 1'b0;
	assign wbs_dat_o = 32'b0;
	assign user_irq = 3'b0;

	eFPGA_top Inst_eFPGA_top(
		.I_top(io_out[37:14]),
		.T_top(io_oeb[37:14]),
		.O_top(io_in[37:14]),
		.A_config_C(),
		.B_config_C(),
		.CLK(io_in[5]),
		.SelfWriteStrobe(1'b0),
		.SelfWriteData(32'b0),
		.Rx(io_in[6]),
		.ComActive(io_out[7]),
		.ReceiveLED(io_out[8]),
		.s_clk(io_in[9]),
		.s_data(io_in[10])
	);
	// unused (shared with caravel)
	assign io_oeb[4:0] = 5'b11111;
	assign io_out[4:0] = 5'b00000;
    // fixed purpose
    assign io_oeb[10:5] = 6'b110011;
    assign io_out[10:9] = 2'b00;
    assign io_out[6:5] = 2'b00;
	// unused currently
	assign io_oeb[13:11] = 3'b111;
	assign io_out[13:11] = 3'b000;

endmodule
